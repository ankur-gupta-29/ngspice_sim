* Simple RC circuit
V1 in 0 PULSE(0 5 0 1n 1n 10n 20n)
R1 in out 1k
C1 out 0 2u
.tran 0.1n 100n
.control
  set filetype=ascii
  run
  write output.raw
  wrdata output.csv time v(out)
  quit
.endc
.end
